
qualquer coisa aqui mesmo
