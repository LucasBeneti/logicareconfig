-- ioweufh
